module moduleName ( ramAddress , ramData );
  

input[15:0] ramAddress;
input[7:0]  ramData;

reg[7:0] firstByte;
reg[7:0] secondByte;

generate
        
endgenerate

generate
        
endgenerate
    
endmodule