module FC(clk,load);
  




    
endmodule